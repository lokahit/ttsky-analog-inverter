magic
tech sky130A
magscale 1 2
timestamp 1756021130
<< error_s >>
rect 2094 1699 2152 1705
rect 2286 1699 2344 1705
rect 2478 1699 2536 1705
rect 2670 1699 2728 1705
rect 2862 1699 2920 1705
rect 3054 1699 3112 1705
rect 3246 1699 3304 1705
rect 3438 1699 3496 1705
rect 3630 1699 3688 1705
rect 3822 1699 3880 1705
rect 2094 1665 2106 1699
rect 2286 1665 2298 1699
rect 2478 1665 2490 1699
rect 2670 1665 2682 1699
rect 2862 1665 2874 1699
rect 3054 1665 3066 1699
rect 3246 1665 3258 1699
rect 3438 1665 3450 1699
rect 3630 1665 3642 1699
rect 3822 1665 3834 1699
rect 2094 1659 2152 1665
rect 2286 1659 2344 1665
rect 2478 1659 2536 1665
rect 2670 1659 2728 1665
rect 2862 1659 2920 1665
rect 3054 1659 3112 1665
rect 3246 1659 3304 1665
rect 3438 1659 3496 1665
rect 3630 1659 3688 1665
rect 3822 1659 3880 1665
rect 1998 1371 2056 1377
rect 2190 1371 2248 1377
rect 2382 1371 2440 1377
rect 2574 1371 2632 1377
rect 2766 1371 2824 1377
rect 2958 1371 3016 1377
rect 3150 1371 3208 1377
rect 3342 1371 3400 1377
rect 3534 1371 3592 1377
rect 3726 1371 3784 1377
rect 1998 1337 2010 1371
rect 2190 1337 2202 1371
rect 2382 1337 2394 1371
rect 2574 1337 2586 1371
rect 2766 1337 2778 1371
rect 2958 1337 2970 1371
rect 3150 1337 3162 1371
rect 3342 1337 3354 1371
rect 3534 1337 3546 1371
rect 3726 1337 3738 1371
rect 1998 1331 2056 1337
rect 2190 1331 2248 1337
rect 2382 1331 2440 1337
rect 2574 1331 2632 1337
rect 2766 1331 2824 1337
rect 2958 1331 3016 1337
rect 3150 1331 3208 1337
rect 3342 1331 3400 1337
rect 3534 1331 3592 1337
rect 3726 1331 3784 1337
rect 2088 459 2146 465
rect 2280 459 2338 465
rect 2472 459 2530 465
rect 2664 459 2722 465
rect 2856 459 2914 465
rect 3048 459 3106 465
rect 3240 459 3298 465
rect 3432 459 3490 465
rect 3624 459 3682 465
rect 3816 459 3874 465
rect 2088 425 2100 459
rect 2280 425 2292 459
rect 2472 425 2484 459
rect 2664 425 2676 459
rect 2856 425 2868 459
rect 3048 425 3060 459
rect 3240 425 3252 459
rect 3432 425 3444 459
rect 3624 425 3636 459
rect 3816 425 3828 459
rect 2088 419 2146 425
rect 2280 419 2338 425
rect 2472 419 2530 425
rect 2664 419 2722 425
rect 2856 419 2914 425
rect 3048 419 3106 425
rect 3240 419 3298 425
rect 3432 419 3490 425
rect 3624 419 3682 425
rect 3816 419 3874 425
rect 1992 149 2050 155
rect 2184 149 2242 155
rect 2376 149 2434 155
rect 2568 149 2626 155
rect 2760 149 2818 155
rect 2952 149 3010 155
rect 3144 149 3202 155
rect 3336 149 3394 155
rect 3528 149 3586 155
rect 3720 149 3778 155
rect 1992 115 2004 149
rect 2184 115 2196 149
rect 2376 115 2388 149
rect 2568 115 2580 149
rect 2760 115 2772 149
rect 2952 115 2964 149
rect 3144 115 3156 149
rect 3336 115 3348 149
rect 3528 115 3540 149
rect 3720 115 3732 149
rect 1992 109 2050 115
rect 2184 109 2242 115
rect 2376 109 2434 115
rect 2568 109 2626 115
rect 2760 109 2818 115
rect 2952 109 3010 115
rect 3144 109 3202 115
rect 3336 109 3394 115
rect 3528 109 3586 115
rect 3720 109 3778 115
<< viali >>
rect 807 1769 905 1824
rect 828 517 925 583
<< metal1 >>
rect 154 1910 4239 2110
rect 394 1617 565 1910
rect 791 1824 918 1910
rect 791 1769 807 1824
rect 905 1769 918 1824
rect 791 1754 918 1769
rect 825 1671 1552 1721
rect 394 1446 823 1617
rect 882 1466 1298 1588
rect 1420 1466 1426 1588
rect 1502 1524 1552 1671
rect 1619 1525 1671 1531
rect 1502 1475 1619 1524
rect 1502 1391 1552 1475
rect 1619 1467 1671 1473
rect 826 1341 1552 1391
rect 258 821 4352 1021
rect 512 374 606 821
rect 810 583 937 821
rect 1680 755 1732 761
rect 1674 703 1680 755
rect 1732 703 1738 755
rect 1680 697 1732 703
rect 810 517 828 583
rect 925 517 937 583
rect 1534 638 1586 644
rect 1534 580 1586 586
rect 810 506 937 517
rect 1535 472 1584 580
rect 848 423 1600 472
rect 512 238 842 374
rect 1298 373 1420 379
rect 907 251 1298 373
rect 1298 245 1420 251
rect 602 197 842 238
rect 1551 162 1600 423
rect 848 113 1600 162
rect 1675 30 1681 82
rect 1733 30 1739 82
rect 1683 -15 1732 30
rect 1641 -174 1773 -15
rect 815 -374 1784 -174
rect 3940 -650 4140 -450
<< via1 >>
rect 1298 1466 1420 1588
rect 1619 1473 1671 1525
rect 1680 703 1732 755
rect 1534 586 1586 638
rect 1298 251 1420 373
rect 1681 30 1733 82
<< metal2 >>
rect 1298 1588 1420 1594
rect 1620 1525 1669 1535
rect 1613 1473 1619 1525
rect 1671 1473 1677 1525
rect 1298 373 1420 1466
rect 1620 1262 1669 1473
rect 1536 1213 1669 1262
rect 1536 753 1585 1213
rect 1680 755 1732 761
rect 1674 753 1680 755
rect 1536 704 1680 753
rect 1536 638 1585 704
rect 1674 703 1680 704
rect 1732 703 1738 755
rect 1680 697 1732 703
rect 1528 586 1534 638
rect 1586 586 1592 638
rect 1292 251 1298 373
rect 1420 251 1426 373
rect 1682 88 1731 697
rect 1681 82 1733 88
rect 1681 24 1733 30
use sky130_fd_pr__pfet_01v8_JBB8V5  XM1
timestamp 1756021130
transform 1 0 856 0 1 1531
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_VL8K8J  XM2
timestamp 1756021130
transform 1 0 878 0 1 292
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_FYAER9  XM3
timestamp 1756021130
transform 1 0 2939 0 1 1518
box -1127 -319 1127 319
use sky130_fd_pr__nfet_01v8_ETUKR2  XM4
timestamp 1756021130
transform 1 0 2933 0 1 287
box -1127 -310 1127 310
<< labels >>
flabel metal1 3940 -650 4140 -450 0 FreeSans 256 0 0 0 output
port 2 nsew
flabel metal1 154 1910 354 2110 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 258 821 458 1021 0 FreeSans 256 0 0 0 VSS
port 1 nsew
flabel metal1 815 -374 1015 -174 0 FreeSans 256 0 0 0 input
port 3 nsew
<< end >>
